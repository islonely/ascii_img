module ascii_img

// fn play_audio(path string) !&ma.Engine {
// 	engine := &ma.Engine{}
// 	result := ma.engine_init(ma.null, engine)
// 	if result != .success {
// 		return error('Failed to initialize audio engine.')
// 	}
// 	if ma.engine_play_sound(engine, path.str, ma.null) != .success {
// 		return error('Failed to load and play "${path}".')
// 	}
// 	ma.engine_uninit(engine)
// }
